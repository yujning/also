// Simple 3-input AND gate test
module test_simple(input a, b, c, output y);
  assign y = a & b & c;
endmodule
